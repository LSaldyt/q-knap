
module us (AL, AZ, AR, CA, CO, CT, DE, FL, GA, ID, IL, IN, IA, KS, KY, LA, ME, MD, MA, MI, MN, MS, MO, MT, NE, NV, NH, NJ, NM, NY, NC, ND, OH, OK, OR, PA, RI, SC, SD, TN, TX, UT, VT, VA, WA, WV, WI, WY, valid);
    input [1:0]AL, AZ, AR, CA, CO, CT, DE, FL, GA, ID, IL, IN, IA, KS, KY, LA, ME, MD, MA, MI, MN, MS, MO, MT, NE, NV, NH, NJ, NM, NY, NC, ND, OH, OK, OR, PA, RI, SC, SD, TN, TX, UT, VT, VA, WA, WV, WI, WY;
    output valid;

    wire [98:0] tests;
    assign tests[0] = WA != OR;
    assign tests[1] = WA != ID;
    assign tests[2] = OR != ID;
    assign tests[3] = OR != CA;
    assign tests[4] = OR != NV;
    assign tests[5] = CA != NV;
    assign tests[6] = CA != AZ;
    assign tests[7] = NV != AZ;
    assign tests[8] = NV != UT;
    assign tests[9] = ID != MT;
    assign tests[10] = ID != WY;
    assign tests[11] = ID != UT;
    assign tests[12] = ID != NV;
    assign tests[13] = UT != WY;
    assign tests[14] = UT != CO;
    assign tests[15] = UT != AZ;
    assign tests[16] = AZ != NM;
    assign tests[17] = MT != WY;
    assign tests[18] = MT != ND;
    assign tests[19] = MT != SD;
    assign tests[20] = WY != SD;
    assign tests[21] = WY != NE;
    assign tests[22] = WY != CO;
    assign tests[23] = CO != KS;
    assign tests[24] = CO != OK;
    assign tests[25] = CO != NM;
    assign tests[26] = NM != OK;
    assign tests[27] = NM != TX;
    assign tests[28] = ND != MN;
    assign tests[29] = ND != SD;
    assign tests[30] = SD != MN;
    assign tests[31] = SD != IA;
    assign tests[32] = SD != NE;
    assign tests[33] = NE != IA;
    assign tests[34] = NE != MO;
    assign tests[35] = NE != KS;
    assign tests[36] = KS != MO;
    assign tests[37] = KS != OK;
    assign tests[38] = OK != MO;
    assign tests[39] = OK != AR;
    assign tests[40] = OK != TX;
    assign tests[41] = TX != AR;
    assign tests[42] = TX != LA;
    assign tests[43] = MN != WI;
    assign tests[44] = MN != IA;
    assign tests[45] = IA != WI;
    assign tests[46] = IA != IL;
    assign tests[47] = IA != MO;
    assign tests[48] = MO != IL;
    assign tests[49] = MO  != KY;
    assign tests[50] = MO != TN;
    assign tests[51] = MO != AR;
    assign tests[52] = AR != MS;
    assign tests[53] = AR != LA;
    assign tests[54] = WI != IL;
    assign tests[55] = WI != MI;
    assign tests[56] = IL != IN;
    assign tests[57] = IL != KY;
    assign tests[58] = MI != IN;
    assign tests[59] = MI != OH;
    assign tests[60] = KY != IN;
    assign tests[61] = KY != OH;
    assign tests[62] = KY != WV;
    assign tests[63] = KY != VA;
    assign tests[64] = KY != TN;
    assign tests[65] = TN != NC;
    assign tests[66] = TN != AL;
    assign tests[67] = TN != MS;
    assign tests[68] = TN != GA;
    assign tests[69] = MS != AL;
    assign tests[70] = AL != GA;
    assign tests[71] = AL != FL;
    assign tests[72] = GA != FL;
    assign tests[73] = SC != GA;
    assign tests[74] = OH != PA;
    assign tests[75] = OH != WV;
    assign tests[76] = WV != OH;
    assign tests[77] = WV != PA;
    assign tests[78] = WV != MD;
    assign tests[79] = WV != VA;
    assign tests[80] = VA != NC;
    assign tests[81] = NC != SC;
    assign tests[82] = PA != MD;
    assign tests[83] = PA != DE;
    assign tests[84] = PA != NJ;
    assign tests[85] = PA != NY;
    assign tests[86] = MD != DE;
    assign tests[87] = DE != NJ;
    assign tests[88] = NJ != NY;
    assign tests[89] = NY != CT;
    assign tests[90] = NY != MA;
    assign tests[91] = NY != VT;
    assign tests[92] = CT != RI;
    assign tests[93] = CT != MA;
    assign tests[94] = VT != NH;
    assign tests[95] = VT != MA;
    assign tests[96] = NH != MA;
    assign tests[97] = NH != ME;
    assign tests[98] = MA != RI;
    assign valid = &tests[98:0];
endmodule
